BZh91AY&SY��B� �_�Py����߰?���P> �  5�5�4d���z�i���昙2h�`��` ���MTd@22 C��  昙2h�`��` ���RD&S&T�T��A�4�dɤ�6`Tv��1�3G��_����B���ܹ�Pc(JT|���f��R{(��cFT��:���m���v^X)z��H��]��uخ�V�~�5�[���f:eL�m��t];pty�
f�eOQ5ƖD0ÕĜzEvIw��թ�;�{�ͨ�%UU�͋���o����a����i0T���'�,��e�H�)�N4��gyU�[�K��������^�j[]t.�y{孳,6����mұfTmB�d/x:��� ��R �I	(��M�ҳ|Z�}lX�l'ΗUf�.�5��_ ��aE��
O�R��0�D!<�%�!�K&�q\$�r7B
��9�~�'=��<7��Sc��|�Tt�����qqx?�������MG�[�K�g'���?�g�wKПB��?i:G��Y�A��x��U
�o����2ǜ���o`�Y�h��4�WR����E&Ř�g5���wMskEI)��7=�&��	RdƓnQ���Y���#�]f��,w��������L%82�MX$���7G�̓|e���L���>��j��b����ýi�x�D����*��pb��F�sa���.��7o��n�$T֨����t�)��){La3�GyR̨�W�^d0NNo7�p�[��%�ƹΞ���f?���(;�X��u��F�7�Ŕ���U�a�,}�y��G��I0e�xkX����J�4r�I����.�a��m�\�ވ�4mqYsq��2w3phc�t�jݺ>����'6��Ҳ5qrX���R��)��RNr�?���)��b8